
//================================================================================================
//    Date         Version  Who  Changes
// -----------------------------------------------------------------------------------------------
// 06-Aug-2022      1.0.0  DWW  Initial creation
//================================================================================================
localparam VERSION_MAJOR = 1;
localparam VERSION_MINOR = 0;
localparam VERSION_BUILD = 0;
localparam VERSION_RCAND = 42;

localparam VERSION_MONTH = 8;
localparam VERSION_DAY   = 6;
localparam VERSION_YEAR  = 2022;
