
`define PBUFF_CHARS         64
`define PBUFF_SIZE          (`PBUFF_CHARS*8)
`define PBUFF_INPUT   input[`PBUFF_SIZE-1:0]
`define PBUFF_OUTPUT output[`PBUFF_SIZE-1:0]
`define PBUFF_REG       reg[`PBUFF_SIZE-1:0]
`define PBUFF_WIRE     wire[`PBUFF_SIZE-1:0]
