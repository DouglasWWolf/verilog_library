
//================================================================================================
//    Date         Version  Who  Changes
// -----------------------------------------------------------------------------------------------
// 27-Jul-2022    1.0.0000  DWW  Initial creation
//================================================================================================
localparam VERSION_MAJOR = 1;
localparam VERSION_MINOR = 0;
localparam VERSION_BUILD = 0;

localparam VERSION_DAY   = 27;
localparam VERSION_MONTH = 7;
localparam VERSION_YEAR  = 2022;
